library verilog;
use verilog.vl_types.all;
entity tb_topall is
end tb_topall;
